// module clint (
//     input               clk,
//     input               rst,

//     input wire[31:0]    inst_i,

//     input reg[63:0]     inst_addr_i, // 用于验证每级传递的pc
//     output reg[63:0]    inst_addr_o, // 用于验证每级传递的pc

//     // from id
//     // input reg[63:0]     csr_raddr_i,
//     input reg[63:0]     csr_waddr_i,
//     input reg[63:0]     csr_data_i,
//     input reg[63:0]     csr_waddr_o,
//     input               csr_wen_o

//     // to ctrl 
//     // output reg[2:0]     stall_flag_o,
//     // output reg[2:0]     flush_flag_o
// );

    


// endmodule