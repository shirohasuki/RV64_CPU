
// module bus_mux (
//     // from IF & MEM
//     input wire      mid_i,
//     input wire[3:0] sid_i,
//     input           wen_i,
//     input           wdata_i,
//     input           waddr_i,
//     input           ren_i,
//     input           raddr_i,

//     // to axi
//     output wire      mid_o,
//     output wire[3:0] sid_o,
//     output           wen_o,
//     output           wdata_o,
//     output           waddr_o,
//     output           ren_o,
//     output           raddr_o,

//     // to IF&MEM
//     output wire[63:0]rdata
// );
// endmodule