// `include "./defines.v"

// module ex_wb(
//     input  wire       clk,
//     input  wire       rst,
    
//     // from ctrl
// //    input  wire       hold_flag_i, // from ctrl 
    
//     //input  wire[31:0] inst_i,    
//     input  wire[63:0] inst_addr_i,    
//     output wire[63:0] inst_addr_o
//     //output wire[31:0] inst_o
// );

//     // dff_set #(32) dff1(clk, rst, 1'b0, `INST_NOP, inst_i, inst_o);

//     dff_set #(64) dff1(clk, rst, 1'b0, 64'b0, inst_addr_i, inst_addr_o);


// endmodule 
