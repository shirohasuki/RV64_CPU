// module id_ram(
//     input  wire       clk,
//     input  wire       rst,

//     // input  wire[31:0] inst_i,       // inst(检测)
//     // input  wire[63:0] inst_addr_i,  // pc(检测)
    
//     output wire[63:0] inst_addr_o,    
//     output wire[31:0] inst_o,
    
//     input wire              mem_wen,
//     input wire[63:0]         mem_waddr_i,
//     input wire              mem_ren,
//     output wire[63:0]        mem_raddr_i 
// );

// 先写成组合
// endmodule