// module uart_tx (
//     input  wire clk,  
//     input  wire rst, 
    
//     input  wire uart_en, 
    
//     output reg txd, 
//     output reg tx_state 
// );

// localparam CLK_Fre = 50_000_000; // 时钟频率
// localparam BAUD = 115200;        // 波特率
// localparam BAUD_DIVISOR = CLK_Fre/BAUD; // 传输一位需要的时钟周期

// always @(posedge clk or negedge rst) begin
    
        
    
// end

// endmodule